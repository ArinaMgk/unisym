// ASCII Verilog Haruno(RFC20)

// 
module shr_ss_byte(
	input A, B,
	output CF, RES);



endmodule
