// ASCII Verilog Haruno(RFC20) [Verilog]

//
module mux_4sel1(// Multiplexer
	input A, B, C, D, SEL0, SEL1,
	output reg RES);
	always @(*)
	begin
		
	end


endmodule
